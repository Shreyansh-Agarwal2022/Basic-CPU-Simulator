//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "new.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w39;    //: /sn:0 {0}(312,568)(330,568)(330,493){1}
//: {2}(330,489)(330,427){3}
//: {4}(330,423)(330,360){5}
//: {6}(330,356)(330,286){7}
//: {8}(330,282)(330,223){9}
//: {10}(330,219)(330,147){11}
//: {12}(330,143)(330,81){13}
//: {14}(330,77)(330,46)(315,46){15}
//: {16}(328,79)(318,79){17}
//: {18}(328,145)(316,145){19}
//: {20}(328,221)(318,221){21}
//: {22}(328,284)(318,284){23}
//: {24}(328,358)(313,358){25}
//: {26}(328,425)(314,425){27}
//: {28}(328,491)(304,491){29}
supply1 w123;    //: /sn:0 {0}(480,1178)(480,1188)(465,1188)(465,1128){1}
reg w101;    //: /sn:0 {0}(-826,471)(-801,471)(-801,518)(-817,518){1}
supply1 w109;    //: /sn:0 {0}(299,1183)(306,1183)(306,1153){1}
supply1 w3;    //: /sn:0 {0}(373,632)(417,632)(417,612){1}
supply0 w19;    //: /sn:0 {0}(-798,672)(-794,672)(-794,695){1}
supply0 w110;    //: /sn:0 {0}(451,1128)(451,1154){1}
supply1 w46;    //: /sn:0 {0}(-466,800)(-440,800){1}
supply0 w67;    //: /sn:0 {0}(-947,344)(-947,341){1}
//: {2}(-947,337)(-947,332){3}
//: {4}(-949,339)(-970,339)(-970,389){5}
//: {6}(-972,391)(-987,391){7}
//: {8}(-970,393)(-970,450)(-939,450)(-939,437){9}
reg w14;    //: /sn:0 {0}(-969,578)(-952,578)(-952,546){1}
supply0 w55;    //: /sn:0 {0}(-234,999)(-215,999)(-215,997){1}
reg w87;    //: /sn:0 {0}(-80,311)(-80,356)(-428,356){1}
//: {2}(-430,354)(-430,299)(-456,299){3}
//: {4}(-430,358)(-430,554)(-328,554){5}
//: {6}(-326,552)(-326,521){7}
//: {8}(-326,556)(-326,557)(-273,557){9}
//: {10}(-269,557)(-214,557)(-214,588)(-187,588){11}
//: {12}(-185,586)(-185,581){13}
//: {14}(-185,590)(-185,631)(-246,631){15}
//: {16}(-248,629)(-248,613){17}
//: {18}(-250,631)(-268,631)(-268,717)(-446,717)(-446,685)(-439,685){19}
//: {20}(-271,555)(-271,548){21}
reg w7;    //: /sn:0 {0}(-116,237)(-110,237)(-110,298)(-96,298){1}
supply0 w117;    //: /sn:0 {0}(-794,785)(-775,785)(-775,805){1}
reg [7:0] w71;    //: /sn:0 {0}(#:-680,522)(-680,532)(-757,532)(-757,567){1}
reg [7:0] w111;    //: /sn:0 {0}(#:367,1183)(367,1206){1}
supply0 w75;    //: /sn:0 {0}(-972,487)(-972,513)(-943,513){1}
supply0 w49;    //: /sn:0 {0}(-817,528)(-801,528)(-801,565){1}
reg [7:0] w47;    //: /sn:0 {0}(#:-995,257)(-995,377){1}
reg [15:0] Instruction16bit;    //: /sn:0 {0}(#:-783,254)(-783,337)(-509,337)(-509,507){1}
//: {2}(-509,508)(-509,534){3}
//: {4}(-509,535)(-509,567){5}
//: {6}(-509,568)(-509,599){7}
//: {8}(-509,600)(-509,630){9}
//: {10}(-509,631)(#:-509,639){11}
wire w16;    //: /sn:0 {0}(362,89)(372,89)(372,104)(327,104)(327,616){1}
wire w58;    //: /sn:0 {0}(-431,816)(-431,857)(-344,857){1}
wire [2:0] w88;    //: /sn:0 {0}(#:-505,568)(-201,568){1}
wire [7:0] w50;    //: /sn:0 {0}(#:-274,971)(-274,985){1}
wire w81;    //: /sn:0 {0}(-323,860)(-44,860){1}
//: {2}(-40,860)(-9,860)(-9,909)(-18,909){3}
//: {4}(-42,862)(-42,910)(-50,910){5}
wire w4;    //: /sn:0 {0}(-978,533)(-962,533){1}
//: {2}(-958,533)(-943,533){3}
//: {4}(-960,531)(-960,370)(-922,370)(-922,278)(-651,278){5}
//: {6}(-647,278)(-96,278){7}
//: {8}(-649,280)(-649,1254)(90,1254)(90,1188)(223,1188){9}
wire [7:0] w56;    //: /sn:0 {0}(#:-140,899)(-140,982){1}
wire w128;    //: /sn:0 {0}(241,1072)(241,1064)(-361,1064)(-361,818){1}
//: {2}(-359,816)(-352,816){3}
//: {4}(-363,816)(-399,816)(-399,826)(-416,826)(-416,816){5}
wire w132;    //: /sn:0 {0}(266,1094)(266,1122)(262,1122)(262,1137){1}
wire w22;    //: /sn:0 {0}(-438,816)(-438,850)(-436,850)(-436,884){1}
//: {2}(-434,886)(-380,886){3}
//: {4}(-436,888)(-436,983)(-309,983)(-309,960){5}
//: {6}(-307,958)(-297,958){7}
//: {8}(-311,958)(-340,958)(-340,1105)(-271,1105){9}
wire w0;    //: /sn:0 {0}(-505,600)(-264,600){1}
wire w20;    //: /sn:0 {0}(312,578)(331,578){1}
wire w29;    //: /sn:0 {0}(318,231)(337,231){1}
wire [2:0] w30;    //: /sn:0 {0}(#:351,645)(351,689)(-148,689)(-148,570){1}
//: {2}(-146,568)(668,568)(#:668,480){3}
//: {4}(-148,566)(-148,558)(#:-172,558){5}
wire w119;    //: /sn:0 {0}(-947,792)(-922,792)(-922,911){1}
wire [7:0] w122;    //: /sn:0 {0}(#:-822,687)(-822,708)(-903,708)(-903,834)(-960,834)(#:-960,808){1}
wire [7:0] w42;    //: /sn:0 {0}(#:279,237)(279,260)(303,260)(303,270)(554,270){1}
//: {2}(558,270)(657,270){3}
//: {4}(556,272)(556,446)(652,446){5}
wire w18;    //: /sn:0 {0}(-380,891)(-442,891)(-442,816){1}
wire w12;    //: /sn:0 {0}(314,435)(362,435){1}
wire w138;    //: /sn:0 {0}(218,1093)(218,1128)(252,1128)(252,1137){1}
wire w54;    //: /sn:0 {0}(-319,977)(-319,999)(-282,999){1}
wire w91;    //: /sn:0 {0}(-423,816)(-423,1065)(-384,1065){1}
wire [2:0] w86;    //: /sn:0 {0}(#:-695,414)(-695,484)(-301,484)(-301,511)(-287,511){1}
wire [7:0] w106;    //: /sn:0 {0}(#:-242,922)(-213,922)(-213,933)(-264,933)(-264,942){1}
wire w31;    //: /sn:0 {0}(318,89)(346,89){1}
wire [7:0] w104;    //: /sn:0 {0}(#:-274,890)(-274,919){1}
//: {2}(-272,921)(-258,921){3}
//: {4}(#:-276,921)(-284,921)(-284,942){5}
wire [7:0] w32;    //: /sn:0 {0}(#:-834,742)(-834,732)(#:-854,732)(-854,641)(-840,641){1}
//: {2}(-838,639)(-838,605)(-854,605){3}
//: {4}(-856,603)(#:-856,534){5}
//: {6}(-858,605)(-892,605){7}
//: {8}(-894,603)(-894,590){9}
//: {10}(-896,605)(-1076,605)(-1076,307)(-1029,307){11}
//: {12}(-1025,307)(#:-965,307){13}
//: {14}(-1027,309)(-1027,377){15}
//: {16}(-838,643)(-838,658){17}
wire [7:0] w68;    //: /sn:0 {0}(#:-146,1210)(-146,1151)(-109,1151)(-109,1122){1}
//: {2}(-107,1120)(-104,1120){3}
//: {4}(-100,1120)(128,1120)(128,778){5}
//: {6}(130,776)(143,776){7}
//: {8}(147,776)(525,776){9}
//: {10}(529,776)(#:739,776)(739,459){11}
//: {12}(#:741,457)(802,457)(802,407){13}
//: {14}(739,455)(739,421){15}
//: {16}(737,457)(#:681,457){17}
//: {18}(527,778)(527,1101)(#:506,1101){19}
//: {20}(145,778)(145,862){21}
//: {22}(126,776)(-53,776){23}
//: {24}(-57,776)(-138,776){25}
//: {26}(-142,776)(-169,776){27}
//: {28}(-171,774)(-171,739){29}
//: {30}(-173,776)(-274,776)(#:-274,874){31}
//: {32}(-140,778)(-140,883){33}
//: {34}(-55,778)(-55,902){35}
//: {36}(-102,1122)(-102,1195)(-142,1195)(-142,1210){37}
//: {38}(-111,1120)(-116,1120){39}
//: {40}(-120,1120)(-131,1120){41}
//: {42}(-135,1120)(-142,1120){43}
//: {44}(-146,1120)(-147,1120){45}
//: {46}(-151,1120)(-153,1120){47}
//: {48}(-157,1120)(-172,1120)(#:-172,1210){49}
//: {50}(-155,1122)(-155,1166)(-169,1166)(-169,1210){51}
//: {52}(-149,1122)(-149,1166)(-165,1166)(-165,1210){53}
//: {54}(-144,1122)(-144,1166)(-161,1166)(-161,1210){55}
//: {56}(-133,1122)(-133,1178)(-154,1178)(-154,1210){57}
//: {58}(-118,1122)(-118,1186)(-150,1186)(-150,1210){59}
wire [7:0] w116;    //: /sn:0 {0}(#:-818,833)(-818,843)(-980,843)(-980,808){1}
wire [7:0] w53;    //: /sn:0 {0}(#:-248,1118)(-248,1189){1}
//: {2}(-246,1191)(-191,1191)(-191,1210){3}
//: {4}(-248,1193)(-248,1201)(-195,1201)(#:-195,1210){5}
wire [7:0] w115;    //: /sn:0 {0}(#:475,1101)(#:490,1101){1}
wire [2:0] w8;    //: /sn:0 {0}(#:-505,535)(-287,535){1}
wire w95;    //: /sn:0 {0}(-235,590)(-218,590)(-218,600)(864,600){1}
wire [2:0] w89;    //: /sn:0 {0}(#:-579,544)(-201,544){1}
wire [7:0] w44;    //: /sn:0 {0}(#:657,264)(462,264)(462,197){1}
//: {2}(464,195)(500,195){3}
//: {4}(504,195)(583,195)(583,440)(#:652,440){5}
//: {6}(502,193)(#:502,183)(501,183)(501,57){7}
//: {8}(460,195)(277,195)(#:277,161){9}
wire w135;    //: /sn:0 {0}(289,1094)(289,1127)(267,1127)(267,1137){1}
wire [7:0] w28;    //: /sn:0 {0}(#:-169,1239)(-169,1280)(-542,1280){1}
//: {2}(-544,1278)(-544,1189){3}
//: {4}(-544,1185)(-544,373)(183,373){5}
//: {6}(185,371)(185,337)(207,337){7}
//: {8}(211,337)(274,337)(#:274,353){9}
//: {10}(209,335)(209,273){11}
//: {12}(211,271)(279,271)(279,279){13}
//: {14}(209,269)(209,202){15}
//: {16}(#:211,200)(279,200)(279,216){17}
//: {18}(209,198)(209,129){19}
//: {20}(#:211,127)(277,127)(277,140){21}
//: {22}(209,125)(209,57)(279,57)(279,74){23}
//: {24}(185,375)(185,410){25}
//: {26}(187,412)(275,412)(#:275,420){27}
//: {28}(185,414)(185,479){29}
//: {30}(#:187,481)(265,481)(265,486){31}
//: {32}(185,483)(#:185,553)(273,553)(273,563){33}
//: {34}(#:-546,1187)(-595,1187)(-595,1171){35}
//: {36}(-546,1280)(-547,1280){37}
wire [7:0] w35;    //: /sn:0 {0}(657,284)(453,284)(#:453,397)(416,397){1}
//: {2}(412,397)(274,397)(#:274,374){3}
//: {4}(414,399)(414,460)(#:652,460){5}
wire [7:0] w45;    //: /sn:0 {0}(#:-885,300)(-885,274){1}
wire w120;    //: /sn:0 {0}(458,1037)(458,1078){1}
wire [7:0] w74;    //: /sn:0 {0}(#:-221,1071)(-199,1071)(-199,1085)(-238,1085)(-238,1089){1}
wire w78;    //: /sn:0 {0}(-404,816)(-404,862)(-344,862){1}
wire [7:0] w2;    //: /sn:0 {0}(#:-180,1210)(-180,1103)(21,1103)(#:21,955){1}
wire [7:0] w41;    //: /sn:0 {0}(#:657,304)(478,304)(478,478){1}
//: {2}(480,480)(#:652,480){3}
//: {4}(478,482)(478,654)(273,654)(#:273,584){5}
wire w11;    //: /sn:0 {0}(378,435)(388,435)(388,450)(361,450)(361,616){1}
wire w129;    //: /sn:0 {0}(243,1093)(243,1122)(257,1122)(257,1137){1}
wire w105;    //: /sn:0 {0}(-1047,361)(-1047,391)(-1035,391){1}
wire [7:0] w83;    //: /sn:0 {0}(#:-922,410)(-888,410){1}
//: {2}(-884,410)(-696,410){3}
//: {4}(-695,410)(-359,410)(-359,488)(-342,488){5}
//: {6}(-886,408)(-886,376){7}
wire w15;    //: /sn:0 {0}(-368,1065)(63,1065)(63,1039){1}
wire w127;    //: /sn:0 {0}(277,882)(277,973){1}
//: {2}(275,975)(270,975){3}
//: {4}(277,977)(277,1028){5}
//: {6}(275,1030)(246,1030)(246,1045){7}
//: {8}(277,1032)(277,1040)(221,1040)(221,1072){9}
wire [7:0] w94;    //: /sn:0 {0}(#:-930,305)(-886,305){1}
//: {2}(-885,305)(-583,305)(-583,543){3}
//: {4}(-583,544)(-583,579){5}
//: {6}(-583,580)(-583,646){7}
//: {8}(-583,647)(-583,663){9}
wire w92;    //: /sn:0 {0}(246,1061)(246,1072){1}
wire [7:0] w43;    //: /sn:0 {0}(#:-970,779)(-970,699)(-1018,699)(-1018,681){1}
//: {2}(-1018,677)(-1018,496)(-856,496)(-856,513){3}
//: {4}(#:-1020,679)(-1093,679)(-1093,652){5}
wire [3:0] w99;    //: /sn:0 {0}(#:-192,1226)(-505,1226)(-505,770)(-418,770){1}
//: {2}(-416,768)(-416,744){3}
//: {4}(#:-414,742)(-337,742)(-337,736){5}
//: {6}(-416,740)(#:-416,698){7}
//: {8}(-416,772)(-416,787){9}
wire [3:0] w100;    //: /sn:0 {0}(#:-579,647)(-406,647)(-406,669){1}
wire w26;    //: /sn:0 {0}(318,294)(344,294){1}
wire [3:0] w76;    //: /sn:0 {0}(#:-505,631)(-426,631)(-426,669){1}
wire w96;    //: /sn:0 {0}(-927,546)(-927,825)(-408,825)(-408,816){1}
wire w125;    //: /sn:0 {0}(458,1021)(458,969){1}
//: {2}(460,967)(485,967)(485,1116)(498,1116)(498,1106){3}
//: {4}(458,965)(458,835)(-397,835)(-397,816){5}
wire w40;    //: /sn:0 {0}(179,869)(191,869)(191,897)(162,897)(162,872){1}
//: {2}(162,868)(162,854)(163,854)(163,847){3}
//: {4}(165,845)(344,845)(344,1032){5}
//: {6}(161,845)(-74,845)(-74,823)(-331,823){7}
//: {8}(160,870)(150,870){9}
wire w6;    //: /sn:0 {0}(304,501)(343,501)(343,500)(359,500){1}
wire [7:0] w13;    //: /sn:0 {0}(#:174,877)(174,991)(#:205,991){1}
wire w114;    //: /sn:0 {0}(-869,767)(-869,785)(-842,785){1}
wire [7:0] w65;    //: /sn:0 {0}(#:-258,1014)(-258,1068){1}
//: {2}(-256,1070)(-237,1070){3}
//: {4}(-258,1072)(-258,1089){5}
wire w34;    //: /sn:0 {0}(260,1158)(260,1178){1}
wire [7:0] w59;    //: /sn:0 {0}(-187,1210)(-187,1089)(-124,1089)(#:-124,1011){1}
wire [7:0] w62;    //: /sn:0 {0}(#:-23,917)(-23,985){1}
wire w25;    //: /sn:0 {0}(360,294)(370,294)(370,309)(347,309)(347,616){1}
wire w72;    //: /sn:0 {0}(-846,672)(-880,672)(-880,655){1}
wire [7:0] w36;    //: /sn:0 {0}(657,277)(445,277)(#:445,327)(405,327){1}
//: {2}(401,327)(279,327)(#:279,300){3}
//: {4}(403,329)(403,453)(#:652,453){5}
wire w82;    //: /sn:0 {0}(-434,816)(-434,877)(-172,877)(-172,866)(-118,866){1}
//: {2}(-114,866)(-86,866)(-86,891)(-103,891){3}
//: {4}(-116,868)(-116,891)(-135,891){5}
wire w124;    //: /sn:0 {0}(264,1073)(264,1042)(-357,1042)(-357,828){1}
//: {2}(-355,826)(-352,826){3}
//: {4}(-359,826)(-393,826)(-393,816){5}
wire w60;    //: /sn:0 {0}(-359,889)(-260,889)(-260,884){1}
//: {2}(-258,882)(-248,882)(-248,889)(-220,889)(-220,880)(-237,880){3}
//: {4}(-262,882)(-269,882){5}
wire [7:0] w112;    //: /sn:0 {0}(-818,817)(#:-818,800){1}
wire w37;    //: /sn:0 {0}(316,155)(343,155){1}
wire [7:0] w73;    //: /sn:0 {0}(#:-176,1210)(-176,1109)(108,1109)(108,1014){1}
//: {2}(108,1010)(108,991)(89,991)(89,975){3}
//: {4}(106,1012)(#:80,1012){5}
wire [7:0] w66;    //: /sn:0 {0}(#:-737,567)(-737,557)(-707,557)(-707,1316)(377,1316)(#:377,1235){1}
wire [7:0] w63;    //: /sn:0 {0}(-184,1210)(-184,1097)(-29,1097)(#:-29,1014){1}
wire w23;    //: /sn:0 {0}(313,368)(338,368){1}
wire w10;    //: /sn:0 {0}(353,231)(363,231)(363,246)(341,246)(341,616){1}
wire [7:0] w70;    //: /sn:0 {0}(#:-802,771)(-802,719)(-747,719)(-747,683){1}
//: {2}(#:-745,681)(-642,681)(-642,665){3}
//: {4}(-747,679)(-747,645){5}
//: {6}(-747,641)(#:-747,596){7}
//: {8}(-749,643)(-806,643)(-806,658){9}
wire [7:0] w84;    //: /sn:0 {0}(#:-1011,406)(-1011,412)(-990,412){1}
//: {2}(-986,412)(-957,412){3}
//: {4}(-988,414)(-988,436)(-1063,436)(-1063,273){5}
wire w24;    //: /sn:0 {0}(-419,816)(-419,853)(-381,853)(-381,821)(-370,821){1}
//: {2}(-366,821)(-352,821){3}
//: {4}(-368,823)(-368,1057)(216,1057)(216,1072){5}
wire w21;    //: /sn:0 {0}(375,500)(385,500)(385,515)(367,515)(367,616){1}
wire [7:0] w108;    //: /sn:0 {0}(#:-834,758)(-834,771){1}
wire w1;    //: /sn:0 {0}(347,578)(374,578)(374,616){1}
wire [7:0] w121;    //: /sn:0 {0}(#:145,878)(145,975)(#:205,975){1}
wire [7:0] w52;    //: /sn:0 {0}(#:-55,918)(-55,985){1}
wire [7:0] w98;    //: /sn:0 {0}(#:686,281)(771,281){1}
//: {2}(775,281)(846,281){3}
//: {4}(850,281)(877,281)(877,584){5}
//: {6}(848,279)(848,242){7}
//: {8}(773,279)(773,263){9}
wire w103;    //: /sn:0 {0}(270,1007)(304,1007){1}
//: {2}(306,1005)(306,928){3}
//: {4}(306,1009)(306,1049)(292,1049)(292,1073){5}
wire w17;    //: /sn:0 {0}(354,368)(386,368)(386,492)(354,492)(354,616){1}
wire w27;    //: /sn:0 {0}(287,1073)(287,1037)(-373,1037)(-373,833){1}
//: {2}(-371,831)(-352,831){3}
//: {4}(-375,831)(-389,831)(-389,816){5}
wire [7:0] w80;    //: /sn:0 {0}(#:-313,498)(897,498)(897,584){1}
wire [7:0] w33;    //: /sn:0 {0}(657,290)(463,290)(#:463,464)(392,464){1}
//: {2}(388,464)(275,464)(#:275,441){3}
//: {4}(390,466)(390,476)(521,476)(521,466)(#:652,466){5}
wire w118;    //: /sn:0 {0}(-401,816)(-401,822)(-394,822)(-394,829){1}
//: {2}(-396,831)(-731,831)(-731,893)(-742,893){3}
//: {4}(-394,833)(-394,1357)(-920,1357)(-920,932){5}
wire w113;    //: /sn:0 {0}(-925,932)(-925,1359)(261,1359)(261,1224){1}
//: {2}(263,1222)(354,1222){3}
//: {4}(261,1220)(261,1199){5}
//: {6}(259,1222)(236,1222)(236,1213)(293,1213){7}
wire w69;    //: /sn:0 {0}(-742,898)(-728,898)(-728,839)(-412,839)(-412,816){1}
wire w48;    //: /sn:0 {0}(-914,523)(-893,523){1}
wire [2:0] w85;    //: /sn:0 {0}(#:-258,525)(673,525)(673,304){1}
wire w90;    //: /sn:0 {0}(26,947)(27,947)(27,932)(-427,932)(-427,816){1}
wire w126;    //: /sn:0 {0}(292,884)(292,989){1}
//: {2}(290,991)(270,991){3}
//: {4}(292,993)(292,1045)(269,1045)(269,1073){5}
wire [7:0] w38;    //: /sn:0 {0}(#:652,433)(596,433)(596,120)(479,120){1}
//: {2}(475,120)(428,120){3}
//: {4}(426,118)(#:426,108)(423,108)(423,51){5}
//: {6}(424,120)(279,120)(#:279,95){7}
//: {8}(477,122)(477,257)(#:657,257){9}
wire [7:0] w5;    //: /sn:0 {0}(657,297)(467,297)(#:467,522)(420,522){1}
//: {2}(418,520)(418,473)(#:652,473){3}
//: {4}(416,522)(265,522)(#:265,507){5}
wire w102;    //: /sn:0 {0}(-67,288)(-23,288){1}
//: {2}(-21,286)(-21,268){3}
//: {4}(-19,266)(4,266){5}
//: {6}(8,266)(16,266)(16,212)(49,212){7}
//: {8}(53,212)(104,212)(104,84)(242,84){9}
//: {10}(51,210)(51,200)(98,200)(98,496)(228,496){11}
//: {12}(51,214)(51,224)(105,224)(105,430)(238,430){13}
//: {14}(6,264)(6,226)(242,226){15}
//: {16}(6,268)(6,280)(21,280)(21,271){17}
//: {18}(23,269)(66,269)(66,573)(236,573){19}
//: {20}(21,267)(21,256)(70,256)(70,150)(240,150){21}
//: {22}(-21,264)(-21,254)(-6,254)(-6,289)(242,289){23}
//: {24}(-21,290)(-21,363)(237,363){25}
wire [7:0] w61;    //: /sn:0 {0}(#:21,939)(21,802){1}
//: {2}(23,800)(40,800){3}
//: {4}(44,800)(172,800){5}
//: {6}(176,800)(385,800){7}
//: {8}(389,800)(410,800){9}
//: {10}(414,800)(#:857,800)(857,647)(887,647)(#:887,613){11}
//: {12}(#:412,802)(412,1103)(440,1103){13}
//: {14}(387,802)(387,1206){15}
//: {16}(174,802)(174,861){17}
//: {18}(42,802)(42,1014)(45,1014){19}
//: {20}(19,800)(-21,800){21}
//: {22}(-25,800)(-79,800){23}
//: {24}(-81,798)(-81,739){25}
//: {26}(-83,800)(-106,800){27}
//: {28}(-110,800)(-242,800)(#:-242,872){29}
//: {30}(-108,802)(-108,883){31}
//: {32}(-23,802)(-23,901){33}
wire [7:0] w64;    //: /sn:0 {0}(#:-49,1014)(-49,1079){1}
//: {2}(-51,1081)(-87,1081)(-87,1075){3}
//: {4}(-49,1083)(-49,1171)(-157,1171)(-157,1210){5}
wire w97;    //: /sn:0 {0}(-579,580)(-264,580){1}
wire w9;    //: /sn:0 {0}(359,155)(369,155)(369,170)(334,170)(334,616){1}
wire w107;    //: /sn:0 {0}(344,1048)(344,1193)(299,1193){1}
wire w79;    //: /sn:0 {0}(-763,895)(-792,895)(-792,583)(-770,583){1}
wire [7:0] w57;    //: /sn:0 {0}(#:-108,899)(-108,982){1}
wire [7:0] w51;    //: /sn:0 {0}(#:-242,888)(-242,985){1}
wire [7:0] w77;    //: /sn:0 {0}(#:-505,508)(-342,508){1}
//: enddecls

  //: LED g116 (w38) @(423,44) /sn:0 /w:[ 5 ] /type:1
  //: LED g164 (w45) @(-885,267) /sn:0 /w:[ 1 ] /type:2
  //: joint g8 (w102) @(-21, 288) /w:[ -1 2 1 24 ]
  _GGREG8 #(10, 10, 20) g4 (.Q(w38), .D(w28), .EN(w31), .CLR(w39), .CK(w102));   //: @(279,84) /sn:0 /w:[ 7 23 0 17 9 ]
  //: GROUND g197 (w117) @(-775,811) /sn:0 /w:[ 1 ]
  assign w97 = w94[3]; //: TAP g157 @(-585,580) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  _GGOR4 #(10) g224 (.I0(w135), .I1(w132), .I2(w129), .I3(w138), .Z(w34));   //: @(260,1148) /sn:0 /R:3 /w:[ 1 1 1 1 0 ]
  //: joint g17 (w28) @(209, 200) /w:[ 16 18 -1 15 ]
  _GGNBUF #(2) g226 (.I(w127), .Z(w92));   //: @(246,1051) /sn:0 /R:3 /w:[ 7 0 ]
  //: joint g137 (w4) @(-649, 278) /w:[ 6 -1 5 8 ]
  //: LED g198 (w114) @(-869,760) /sn:0 /w:[ 0 ] /type:0
  _GGNBUF8 #(2) g92 (.I(w65), .Z(w74));   //: @(-231,1071) /sn:0 /w:[ 3 0 ]
  _GGBUFIF8 #(4, 6) g74 (.Z(w56), .I(w68), .E(w82));   //: @(-140,889) /sn:0 /R:3 /w:[ 0 33 5 ]
  //: joint g30 (w39) @(330, 221) /w:[ -1 10 20 9 ]
  //: joint g183 (w98) @(848, 281) /w:[ 4 6 3 -1 ]
  _GGROM8x8 #(10, 30) g130 (.A(w32), .D(w94), .OE(w67));   //: @(-947,306) /sn:0 /w:[ 13 0 3 ] /mem:"/home/linux/Downloads/instruction.mem"
  //: joint g77 (w68) @(-140, 776) /w:[ 25 -1 26 32 ]
  _GGREG8 #(10, 10, 20) g1 (.Q(w42), .D(w28), .EN(w29), .CLR(w39), .CK(w102));   //: @(279,226) /sn:0 /w:[ 0 17 0 21 15 ]
  Comp g111 (.a(w121), .b(w13), .et(w127), .gt(w126), .lt(w103));   //: @(206, 959) /sz:(63, 64) /sn:0 /p:[ Li0>1 Li1>1 Ro0<3 Ro1<3 Ro2<0 ]
  //: joint g214 (w61) @(412, 800) /w:[ 10 -1 9 12 ]
  //: joint g179 (w68) @(-171, 776) /w:[ 27 28 30 -1 ]
  //: joint g144 (w87) @(-248, 631) /w:[ 15 16 18 -1 ]
  _GGNBUF #(2) g51 (.I(w17), .Z(w23));   //: @(348,368) /sn:0 /R:2 /w:[ 0 1 ]
  //: joint g190 (w68) @(-102, 1120) /w:[ 4 -1 3 36 ]
  //: joint g206 (w118) @(-394, 831) /w:[ -1 1 2 4 ]
  //: SWITCH g161 (w7) @(-133,237) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g70 (w54) @(-319,970) /sn:0 /w:[ 0 ] /type:0
  _GGROM8x8 #(10, 30) g149 (.A(w84), .D(w83), .OE(w67));   //: @(-939,411) /sn:0 /w:[ 3 0 9 ] /mem:"/home/linux/Downloads/instruction.mem"
  _GGBUFIF8 #(4, 6) g65 (.Z(w104), .I(w68), .E(w60));   //: @(-274,880) /sn:0 /R:3 /w:[ 0 31 5 ]
  //: joint g25 (w39) @(330, 79) /w:[ -1 14 16 13 ]
  //: joint g10 (w102) @(51, 212) /w:[ 8 10 7 12 ]
  _GGBUFIF8 #(4, 6) g103 (.Z(w13), .I(w61), .E(w40));   //: @(174,867) /sn:0 /R:3 /w:[ 0 17 0 ]
  //: joint g220 (w125) @(458, 967) /w:[ 2 4 -1 1 ]
  assign w76 = Instruction16bit[15:12]; //: TAP g64 @(-511,631) /sn:0 /R:2 /w:[ 0 10 9 ] /ss:1
  _GGMUX2x8 #(8, 8) g185 (.I0(w111), .I1(w61), .S(w113), .Z(w66));   //: @(377,1222) /sn:0 /w:[ 1 15 3 1 ] /ss:0 /do:0
  _GGNBUF #(2) g49 (.I(w9), .Z(w37));   //: @(353,155) /sn:0 /R:2 /w:[ 0 1 ]
  _GGDECODER15 #(6, 6) g72 (.I(w99), .E(w46), .Z0(w18), .Z1(w22), .Z2(w82), .Z3(w58), .Z4(w90), .Z5(w91), .Z6(w24), .Z7(w128), .Z8(w69), .Z9(w96), .Z10(w78), .Z11(w118), .Z12(w125), .Z13(w124), .Z14(w27));   //: @(-416,800) /sn:0 /w:[ 9 1 1 0 0 0 1 0 0 5 1 1 0 0 5 5 5 ] /ss:0 /do:0
  //: joint g136 (w81) @(-42, 860) /w:[ 2 -1 1 4 ]
  _GGMUX2 #(8, 8) g142 (.I0(w0), .I1(w97), .S(w87), .Z(w95));   //: @(-248,590) /sn:0 /R:1 /w:[ 1 1 17 0 ] /ss:0 /do:0
  _GGREG8 #(10, 10, 20) g6 (.Q(w5), .D(w28), .EN(w6), .CLR(w39), .CK(w102));   //: @(265,496) /sn:0 /w:[ 5 31 0 29 11 ]
  _GGMUX2x8 #(8, 8) g124 (.I0(w71), .I1(w66), .S(w79), .Z(w70));   //: @(-747,583) /sn:0 /w:[ 1 0 1 7 ] /ss:0 /do:0
  //: joint g35 (w44) @(462, 195) /w:[ 2 -1 8 1 ]
  _GGREG8 #(10, 10, 20) g7 (.Q(w41), .D(w28), .EN(w20), .CLR(w39), .CK(w102));   //: @(273,573) /sn:0 /w:[ 5 33 0 0 19 ]
  assign w0 = Instruction16bit[11]; //: TAP g58 @(-511,600) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: joint g229 (w103) @(306, 1007) /w:[ -1 2 1 4 ]
  //: joint g200 (w68) @(-133, 1120) /w:[ 41 -1 42 56 ]
  //: joint g181 (w61) @(-81, 800) /w:[ 23 24 26 -1 ]
  //: LED g98 (w73) @(89,968) /sn:0 /w:[ 3 ] /type:1
  //: LED g192 (w44) @(501,50) /sn:0 /w:[ 7 ] /type:1
  //: joint g204 (w70) @(-747, 643) /w:[ -1 6 8 5 ]
  //: LED g85 (w64) @(-87,1068) /sn:0 /w:[ 3 ] /type:3
  //: joint g67 (w60) @(-260, 882) /w:[ 2 -1 4 1 ]
  //: GROUND g126 (w19) @(-794,701) /sn:0 /w:[ 1 ]
  //: joint g208 (w43) @(-1018, 679) /w:[ -1 2 4 1 ]
  _GGNBUF #(2) g54 (.I(w1), .Z(w20));   //: @(341,578) /sn:0 /R:2 /w:[ 0 1 ]
  //: joint g33 (w38) @(477, 120) /w:[ 1 -1 2 8 ]
  _GGBUFIF8 #(4, 6) g81 (.Z(w62), .I(w61), .E(w81));   //: @(-23,907) /sn:0 /R:3 /w:[ 0 33 3 ]
  _GGNBUF #(2) g52 (.I(w11), .Z(w12));   //: @(372,435) /sn:0 /R:2 /w:[ 0 1 ]
  //: joint g40 (w42) @(556, 270) /w:[ 2 -1 1 4 ]
  //: joint g163 (w87) @(-430, 356) /w:[ 1 2 -1 4 ]
  //: frame g132 @(-1161,214) /sn:0 /wi:672 /ht:507 /tx:"Program Counter"
  _GGAND2 #(6) g222 (.I0(w103), .I1(w27), .Z(w135));   //: @(289,1084) /sn:0 /R:3 /w:[ 5 0 0 ]
  //: GROUND g217 (w110) @(451,1160) /sn:0 /w:[ 1 ]
  //: joint g210 (w70) @(-747, 681) /w:[ 2 4 -1 1 ]
  //: joint g12 (w102) @(-21, 266) /w:[ 4 22 -1 3 ]
  //: joint g108 (w61) @(174, 800) /w:[ 6 -1 5 16 ]
  //: GROUND g131 (w67) @(-947,350) /sn:0 /w:[ 0 ]
  //: joint g106 (w40) @(162, 870) /w:[ -1 2 8 1 ]
  //: joint g230 (w24) @(-368, 821) /w:[ 2 -1 1 4 ]
  _GGADD8 #(68, 70, 62, 64) g194 (.A(w108), .B(w70), .S(w112), .CI(w117), .CO(w114));   //: @(-818,787) /sn:0 /w:[ 1 0 1 0 1 ]
  //: SWITCH g177 (w14) @(-986,578) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g228 (w126) @(292, 991) /w:[ -1 1 2 4 ]
  //: LED g209 (w70) @(-642,658) /sn:0 /w:[ 3 ] /type:3
  _GGROM8x8 #(10, 30) g96 (.A(w61), .D(w73), .OE(w15));   //: @(63,1013) /sn:0 /w:[ 19 5 1 ] /mem:"/home/linux/Downloads/memory.mem"
  //: joint g221 (w44) @(502, 195) /w:[ 4 6 3 -1 ]
  //: LED g114 (w126) @(292,877) /sn:0 /w:[ 0 ] /type:0
  _GGNBUF8 #(2) g196 (.I(w32), .Z(w108));   //: @(-834,748) /sn:0 /R:3 /w:[ 0 0 ]
  //: joint g19 (w28) @(185, 412) /w:[ 26 25 -1 28 ]
  //: joint g117 (w68) @(-144, 1120) /w:[ 43 -1 44 54 ]
  //: joint g78 (w61) @(-108, 800) /w:[ 27 -1 28 30 ]
  //: LED g125 (w72) @(-880,648) /sn:0 /w:[ 1 ] /type:0
  _GGAND2 #(6) g223 (.I0(w127), .I1(w24), .Z(w138));   //: @(218,1083) /sn:0 /R:3 /w:[ 9 5 0 ]
  //: joint g113 (w68) @(-109, 1120) /w:[ 2 -1 38 1 ]
  //: joint g219 (w68) @(-118, 1120) /w:[ 39 -1 40 58 ]
  //: joint g63 (w98) @(773, 281) /w:[ 2 8 1 -1 ]
  assign w100 = w94[7:4]; //: TAP g155 @(-585,647) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  _GGNBUF #(2) g100 (.I(w91), .Z(w15));   //: @(-378,1065) /sn:0 /w:[ 1 0 ]
  //: joint g93 (w99) @(-416, 770) /w:[ -1 2 1 8 ]
  _GGOR4 #(10) g105 (.I0(w128), .I1(w24), .I2(w124), .I3(w27), .Z(w40));   //: @(-341,823) /sn:0 /w:[ 3 3 3 3 7 ]
  _GGBUFIF8 #(4, 6) g215 (.Z(w115), .I(w68), .E(w125));   //: @(500,1101) /sn:0 /R:2 /w:[ 1 19 3 ]
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g212 (.A(w61), .D(w115), .WE(w120), .OE(w123), .CS(w110));   //: @(458,1102) /sn:0 /w:[ 13 0 1 1 0 ]
  //: joint g211 (w4) @(-960, 533) /w:[ 2 4 1 -1 ]
  //: LED g205 (w113) @(300,1213) /sn:0 /R:3 /w:[ 7 ] /type:0
  //: joint g38 (w68) @(739, 457) /w:[ 12 14 16 11 ]
  _GGBUFIF8 #(4, 6) g101 (.Z(w2), .I(w61), .E(w90));   //: @(21,945) /sn:0 /R:3 /w:[ 1 0 0 ]
  //: joint g43 (w35) @(414, 397) /w:[ 1 -1 2 4 ]
  _GGREG8 #(10, 10, 20) g0 (.Q(w44), .D(w28), .EN(w37), .CLR(w39), .CK(w102));   //: @(277,150) /sn:0 /w:[ 9 21 0 19 21 ]
  //: joint g48 (w39) @(330, 491) /w:[ -1 2 28 1 ]
  //: frame g37 @(17,1) /sn:0 /wi:929 /ht:713 /tx:"Register File"
  _GGCLOCK_P10000_0_50 g122 (.Z(w4));   //: @(-991,533) /sn:0 /w:[ 0 ] /omega:10000 /phi:0 /duty:50
  //: GROUND g120 (w49) @(-801,571) /sn:0 /w:[ 1 ]
  _GGBUFIF8 #(4, 6) g80 (.Z(w52), .I(w68), .E(w81));   //: @(-55,908) /sn:0 /R:3 /w:[ 0 35 5 ]
  //: joint g95 (w28) @(185, 373) /w:[ -1 6 5 24 ]
  //: joint g76 (w82) @(-116, 866) /w:[ 2 -1 1 4 ]
  _GGNBUF #(2) g189 (.I(w40), .Z(w107));   //: @(344,1038) /sn:0 /R:3 /w:[ 5 0 ]
  //: LED g178 (w68) @(-171,732) /sn:0 /w:[ 29 ] /type:3
  //: joint g170 (w84) @(-988, 412) /w:[ 2 -1 1 4 ]
  //: LED g152 (w105) @(-1047,354) /sn:0 /w:[ 0 ] /type:0
  _GGBUFIF8 #(4, 6) g75 (.Z(w57), .I(w61), .E(w82));   //: @(-108,889) /sn:0 /R:3 /w:[ 0 31 3 ]
  //: joint g44 (w33) @(390, 464) /w:[ 1 -1 2 4 ]
  //: LED g182 (w98) @(848,235) /sn:0 /w:[ 7 ] /type:1
  assign w86 = w83[7:5]; //: TAP g159 @(-695,408) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g47 (w39) @(330, 425) /w:[ -1 4 26 3 ]
  //: joint g16 (w28) @(209, 127) /w:[ 20 22 -1 19 ]
  _GGREG8 #(10, 10, 20) g3 (.Q(w35), .D(w28), .EN(w23), .CLR(w39), .CK(w102));   //: @(274,363) /sn:0 /w:[ 3 9 0 25 25 ]
  _GGMUX2x4 #(8, 8) g143 (.I0(w76), .I1(w100), .S(w87), .Z(w99));   //: @(-416,685) /sn:0 /w:[ 1 1 19 7 ] /ss:0 /do:0
  //: DIP Default2 (w71) @(-680,512) /sn:0 /w:[ 0 ] /st:2 /dn:1
  _GGDECODER8 #(6, 6) g26 (.I(w30), .E(w3), .Z0(w1), .Z1(w21), .Z2(w11), .Z3(w17), .Z4(w25), .Z5(w10), .Z6(w9), .Z7(w16));   //: @(351,632) /sn:0 /R:2 /w:[ 0 0 1 1 1 1 1 1 1 1 ] /ss:0 /do:0
  //: joint g109 (w68) @(128, 776) /w:[ 6 -1 22 5 ]
  //: joint g90 (w32) @(-856, 605) /w:[ 3 4 6 -1 ]
  //: joint g174 (w28) @(-544, 1187) /w:[ -1 4 34 3 ]
  //: joint g158 (w67) @(-970, 391) /w:[ -1 5 6 8 ]
  //: joint g128 (w32) @(-894, 605) /w:[ 7 8 10 -1 ]
  _GGREG8 #(10, 10, 20) g2 (.Q(w36), .D(w28), .EN(w26), .CLR(w39), .CK(w102));   //: @(279,289) /sn:0 /w:[ 3 13 0 23 23 ]
  _GGNBUF #(2) g23 (.I(w16), .Z(w31));   //: @(356,89) /sn:0 /R:2 /w:[ 0 1 ]
  _GGMUX15x8 #(34, 34) g91 (.I0(w53), .I1(w53), .I2(w59), .I3(w63), .I4(w2), .I5(w73), .I6(w68), .I7(w68), .I8(w68), .I9(w68), .I10(w64), .I11(w68), .I12(w68), .I13(w68), .I14(w68), .S(w99), .Z(w28));   //: @(-169,1226) /sn:0 /w:[ 5 3 0 0 0 0 49 51 53 55 5 57 59 0 37 0 0 ] /ss:0 /do:0
  _GGMUX2x8 #(8, 8) g127 (.I0(w65), .I1(w74), .S(w22), .Z(w53));   //: @(-248,1105) /sn:0 /w:[ 5 1 9 0 ] /ss:0 /do:0
  _GGMUX2x3 #(8, 8) g141 (.I0(w88), .I1(w89), .S(w87), .Z(w30));   //: @(-185,558) /sn:0 /R:1 /w:[ 1 1 13 5 ] /ss:0 /do:0
  _GGMUX2x8 #(8, 8) g86 (.I0(w98), .I1(w80), .S(w95), .Z(w61));   //: @(887,600) /sn:0 /w:[ 5 1 1 11 ] /ss:0 /do:0
  //: SWITCH g24 (w39) @(298,46) /sn:0 /w:[ 15 ] /st:1 /dn:1
  //: VDD g39 (w3) @(428,612) /sn:0 /w:[ 1 ]
  _GGBUFIF8 #(4, 6) g104 (.Z(w121), .I(w68), .E(w40));   //: @(145,868) /sn:0 /R:3 /w:[ 0 21 9 ]
  assign w77 = Instruction16bit[7:0]; //: TAP g60 @(-511,508) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: joint g110 (w68) @(-155, 1120) /w:[ 47 -1 48 50 ]
  //: LED g121 (w43) @(-1093,645) /sn:0 /w:[ 5 ] /type:3
  //: joint g29 (w39) @(330, 145) /w:[ -1 12 18 11 ]
  //: joint g168 (w67) @(-947, 339) /w:[ -1 2 4 1 ]
  //: joint g18 (w28) @(209, 337) /w:[ 8 10 7 -1 ]
  _GGOR2 #(6) g82 (.I0(w58), .I1(w78), .Z(w81));   //: @(-333,860) /sn:0 /w:[ 1 1 0 ]
  //: joint g199 (w113) @(261, 1222) /w:[ 2 4 6 1 ]
  //: joint g94 (w28) @(-544, 1280) /w:[ 1 2 36 -1 ]
  _GGREG8 #(10, 10, 20) g119 (.Q(w32), .D(w43), .EN(w49), .CLR(w101), .CK(w48));   //: @(-856,523) /sn:0 /w:[ 5 3 0 1 1 ]
  //: joint g173 (w104) @(-274, 921) /w:[ 2 1 4 -1 ]
  //: joint g154 (w53) @(-248, 1191) /w:[ 2 1 -1 4 ]
  //: LED g166 (w83) @(-886,369) /sn:0 /w:[ 7 ] /type:2
  //: joint g107 (w68) @(145, 776) /w:[ 8 -1 7 20 ]
  _GGNBUF8 #(2) g172 (.I(w104), .Z(w106));   //: @(-252,922) /sn:0 /w:[ 3 0 ]
  //: LED g184 (w68) @(802,400) /sn:0 /w:[ 13 ] /type:1
  //: joint g188 (w40) @(163, 845) /w:[ 4 -1 6 3 ]
  //: joint g216 (w68) @(527, 776) /w:[ 10 -1 9 18 ]
  _GGAND2 #(6) g193 (.I0(w126), .I1(w124), .Z(w132));   //: @(266,1084) /sn:0 /R:3 /w:[ 5 0 0 ]
  _GGNBUF #(2) g50 (.I(w25), .Z(w26));   //: @(354,294) /sn:0 /R:2 /w:[ 0 1 ]
  //: joint g68 (w22) @(-309, 958) /w:[ 6 -1 8 5 ]
  _GGMUX2 #(8, 8) g133 (.I0(w4), .I1(w75), .S(w96), .Z(w48));   //: @(-927,523) /sn:0 /R:1 /w:[ 3 1 0 0 ] /ss:0 /do:0
  _GGMUL8 #(124) g73 (.A(w56), .B(w57), .P(w59));   //: @(-124,998) /sn:0 /w:[ 1 1 1 ]
  //: joint g9 (w102) @(6, 266) /w:[ 6 14 5 16 ]
  //: joint g225 (w127) @(277, 975) /w:[ -1 1 2 4 ]
  _GGAND2 #(6) g102 (.I0(w92), .I1(w128), .Z(w129));   //: @(243,1083) /sn:0 /R:3 /w:[ 1 0 0 ]
  //: joint g186 (w61) @(387, 800) /w:[ 8 -1 7 14 ]
  //: LED g169 (w84) @(-1063,266) /sn:0 /w:[ 5 ] /type:1
  _GGOR2 #(6) g71 (.I0(w22), .I1(w18), .Z(w60));   //: @(-369,889) /sn:0 /w:[ 3 0 0 ]
  _GGNBUF #(2) g22 (.I(w10), .Z(w29));   //: @(347,231) /sn:0 /R:2 /w:[ 0 1 ]
  //: joint g31 (w39) @(330, 284) /w:[ -1 8 22 7 ]
  assign w8 = Instruction16bit[7:5]; //: TAP g59 @(-511,535) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g231 (w128) @(-361, 816) /w:[ 2 -1 4 1 ]
  //: DIP g87 (w111) @(367,1173) /sn:0 /w:[ 0 ] /st:2 /dn:1
  //: LED g180 (w61) @(-81,732) /sn:0 /w:[ 25 ] /type:3
  //: joint g99 (w73) @(108, 1012) /w:[ -1 2 4 1 ]
  //: joint g83 (w68) @(-55, 776) /w:[ 23 -1 24 34 ]
  //: joint g203 (w32) @(-838, 641) /w:[ -1 2 1 16 ]
  //: LED g36 (w68) @(739,414) /sn:0 /w:[ 15 ] /type:3
  //: joint g45 (w5) @(418, 522) /w:[ 1 2 4 -1 ]
  _GGMUX8x8 #(20, 20) g41 (.I0(w41), .I1(w5), .I2(w33), .I3(w35), .I4(w36), .I5(w42), .I6(w44), .I7(w38), .S(w30), .Z(w68));   //: @(668,457) /sn:0 /R:1 /w:[ 3 3 5 5 5 5 5 0 3 17 ] /ss:0 /do:0
  _GGREG #(10, 10, 20) g138 (.Q(w113), .D(w34), .EN(w107), .CLR(w109), .CK(w4));   //: @(260,1188) /sn:0 /w:[ 5 1 1 0 9 ]
  //: LED g69 (w28) @(-595,1164) /sn:0 /w:[ 35 ] /type:3
  //: joint g42 (w36) @(403, 327) /w:[ 1 -1 2 4 ]
  assign w89 = w94[2:0]; //: TAP g156 @(-585,544) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  _GGNBUF #(2) g213 (.I(w125), .Z(w120));   //: @(458,1027) /sn:0 /R:3 /w:[ 0 0 ]
  //: joint g151 (w32) @(-1027, 307) /w:[ 12 -1 11 14 ]
  _GGBUFIF8 #(4, 6) g66 (.Z(w51), .I(w61), .E(w60));   //: @(-242,878) /sn:0 /R:3 /w:[ 0 29 3 ]
  //: joint g167 (w83) @(-886, 410) /w:[ 2 6 1 -1 ]
  //: joint g233 (w27) @(-373, 831) /w:[ 2 -1 4 1 ]
  //: joint g232 (w124) @(-357, 826) /w:[ 2 -1 4 1 ]
  //: joint g191 (w38) @(426, 120) /w:[ 3 4 6 -1 ]
  _GGMUX2 #(8, 8) g162 (.I0(w7), .I1(w4), .S(w87), .Z(w102));   //: @(-80,288) /sn:0 /R:1 /w:[ 1 7 0 0 ] /ss:0 /do:0
  //: joint g146 (w87) @(-271, 557) /w:[ 10 20 9 -1 ]
  //: joint g153 (w65) @(-258, 1070) /w:[ 2 1 -1 4 ]
  //: GROUND g57 (w55) @(-215,991) /sn:0 /R:2 /w:[ 1 ]
  _GGADD8 #(68, 70, 62, 64) g34 (.A(w50), .B(w51), .S(w65), .CI(w55), .CO(w54));   //: @(-258,1001) /sn:0 /w:[ 1 1 0 0 1 ]
  //: VDD g28 (w46) @(-466,789) /sn:0 /R:1 /w:[ 0 ]
  //: joint g46 (w41) @(478, 480) /w:[ 2 1 -1 4 ]
  _GGADD8 #(68, 70, 62, 64) g150 (.A(w32), .B(w47), .S(w84), .CI(w67), .CO(w105));   //: @(-1011,393) /sn:0 /w:[ 15 1 0 7 1 ]
  //: frame g118 @(-522,765) /sn:0 /wi:1081 /ht:506 /tx:"ALU"
  //: joint g84 (w61) @(-23, 800) /w:[ 21 -1 22 32 ]
  //: joint g11 (w102) @(21, 269) /w:[ 18 20 -1 17 ]
  _GGREG8 #(10, 10, 20) g5 (.Q(w33), .D(w28), .EN(w12), .CLR(w39), .CK(w102));   //: @(275,430) /sn:0 /w:[ 3 27 0 27 13 ]
  //: joint g14 (w61) @(21, 800) /w:[ 2 -1 20 1 ]
  _GGAND2 #(6) g201 (.I0(w113), .I1(w118), .Z(w119));   //: @(-922,921) /sn:0 /R:1 /w:[ 0 5 1 ]
  //: LED g112 (w103) @(306,921) /sn:0 /w:[ 3 ] /type:0
  //: VDD g187 (w109) @(317,1153) /sn:0 /w:[ 1 ]
  //: LED g61 (w98) @(773,256) /sn:0 /w:[ 9 ] /type:3
  //: LED g123 (w32) @(-894,583) /sn:0 /w:[ 9 ] /type:1
  _GGMUX8x8 #(20, 20) g21 (.I0(w41), .I1(w5), .I2(w33), .I3(w35), .I4(w36), .I5(w42), .I6(w44), .I7(w38), .S(w85), .Z(w98));   //: @(673,281) /sn:0 /R:1 /w:[ 0 0 0 0 0 3 0 9 1 0 ] /ss:0 /do:0
  //: LED g115 (w127) @(277,875) /sn:0 /w:[ 0 ] /type:0
  //: joint g20 (w28) @(185, 481) /w:[ 30 29 -1 32 ]
  //: joint g32 (w39) @(330, 358) /w:[ -1 6 24 5 ]
  _GGDIV8 #(236, 236) g79 (.A(w52), .B(w62), .Q(w63), .R(w64));   //: @(-39,1001) /sn:0 /w:[ 1 1 1 0 ]
  //: joint g176 (w99) @(-416, 742) /w:[ 4 6 -1 3 ]
  //: LED g175 (w99) @(-337,729) /sn:0 /w:[ 5 ] /type:1
  //: joint g97 (w61) @(42, 800) /w:[ 4 -1 3 18 ]
  //: GROUND g134 (w75) @(-972,481) /sn:0 /R:2 /w:[ 0 ]
  //: joint g145 (w87) @(-185, 588) /w:[ -1 12 11 14 ]
  //: DIP g129 (w47) @(-995,247) /sn:0 /w:[ 0 ] /st:1 /dn:1
  _GGADD8 #(68, 70, 62, 64) g89 (.A(w32), .B(w70), .S(w122), .CI(w19), .CO(w72));   //: @(-822,674) /sn:0 /w:[ 17 9 0 0 0 ]
  //: joint g15 (w28) @(209, 271) /w:[ 12 14 -1 11 ]
  //: SWITCH g148 (w87) @(-473,299) /sn:0 /w:[ 3 ] /st:1 /dn:1
  //: joint g227 (w127) @(277, 1030) /w:[ -1 5 6 8 ]
  _GGMUX2x8 #(8, 8) g202 (.I0(w122), .I1(w116), .S(w119), .Z(w43));   //: @(-970,792) /sn:0 /R:2 /w:[ 1 1 0 0 ] /ss:0 /do:0
  assign w45 = w94[7:0]; //: TAP g165 @(-885,303) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  //: joint g147 (w87) @(-326, 554) /w:[ -1 6 5 8 ]
  //: joint g27 (w22) @(-436, 886) /w:[ 2 1 -1 4 ]
  //: SWITCH g160 (w101) @(-843,471) /sn:0 /w:[ 0 ] /st:1 /dn:1
  assign w88 = Instruction16bit[10:8]; //: TAP g62 @(-511,568) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  _GGMUX2x8 #(8, 8) g171 (.I0(w104), .I1(w106), .S(w22), .Z(w50));   //: @(-274,958) /sn:0 /w:[ 5 1 7 0 ] /ss:0 /do:0
  //: VDD g218 (w123) @(491,1178) /sn:0 /w:[ 0 ]
  _GGNBUF8 #(2) g195 (.I(w112), .Z(w116));   //: @(-818,823) /sn:0 /R:3 /w:[ 0 0 ]
  //: DIP g55 (Instruction16bit) @(-783,244) /sn:0 /w:[ 0 ] /st:51457 /dn:1
  //: joint g88 (w68) @(-149, 1120) /w:[ 45 -1 46 52 ]
  //: joint g135 (w64) @(-49, 1081) /w:[ -1 1 2 4 ]
  _GGNBUF #(2) g53 (.I(w21), .Z(w6));   //: @(369,500) /sn:0 /R:2 /w:[ 0 1 ]
  //: joint g13 (w30) @(-148, 568) /w:[ 2 4 -1 1 ]
  _GGMUX2x8 #(8, 8) g139 (.I0(w77), .I1(w83), .S(w87), .Z(w80));   //: @(-326,498) /sn:0 /R:1 /w:[ 1 5 7 0 ] /ss:0 /do:0
  _GGMUX2x3 #(8, 8) g140 (.I0(w8), .I1(w86), .S(w87), .Z(w85));   //: @(-271,525) /sn:0 /R:1 /w:[ 1 1 21 0 ] /ss:0 /do:0
  _GGOR2 #(6) g207 (.I0(w69), .I1(w118), .Z(w79));   //: @(-753,895) /sn:0 /R:2 /w:[ 0 3 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin comp4
module comp4(b1, b2, g, b3, a1, l, e, a0, a2, a3, b0);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input a2;    //: /sn:0 {0}(75,-51)(152,-51){1}
//: {2}(156,-51)(178,-51){3}
//: {4}(154,-49)(154,-3)(236,-3){5}
input b2;    //: /sn:0 {0}(77,2)(143,2){1}
//: {2}(147,2)(178,2){3}
//: {4}(145,0)(145,-46)(236,-46){5}
input a3;    //: /sn:0 {0}(74,-155)(149,-155){1}
//: {2}(153,-155)(178,-155){3}
//: {4}(151,-153)(151,-112)(235,-112){5}
output l;    //: /sn:0 {0}(604,28)(571,28)(571,28)(664,28){1}
input b3;    //: /sn:0 {0}(73,-107)(141,-107){1}
//: {2}(145,-107)(178,-107){3}
//: {4}(143,-109)(143,-150)(236,-150){5}
input a1;    //: /sn:0 {0}(80,57)(154,57){1}
//: {2}(158,57)(178,57){3}
//: {4}(156,59)(156,106)(236,106){5}
input b1;    //: /sn:0 {0}(80,111)(145,111){1}
//: {2}(149,111)(178,111){3}
//: {4}(147,109)(147,62)(236,62){5}
input a0;    //: /sn:0 {0}(236,207)(158,207)(158,158){1}
//: {2}(160,156)(178,156){3}
//: {4}(156,156)(81,156){5}
input b0;    //: /sn:0 {0}(83,212)(146,212){1}
//: {2}(150,212)(178,212){3}
//: {4}(148,210)(148,161)(236,161){5}
output e;    //: /sn:0 {0}(449,268)(631,268)(631,268)(669,268){1}
output g;    //: /sn:0 {0}(601,172)(620,172)(620,172)(666,172){1}
wire w16;    //: /sn:0 {0}(257,-48)(306,-48){1}
//: {2}(308,-50)(308,-88)(428,-88){3}
//: {4}(308,-46)(308,-29)(323,-29){5}
wire w6;    //: /sn:0 {0}(428,266)(380,266)(380,212){1}
//: {2}(382,210)(428,210){3}
//: {4}(380,208)(380,158){5}
//: {6}(382,156)(428,156){7}
//: {8}(380,154)(380,104){9}
//: {10}(382,102)(428,102){11}
//: {12}(380,100)(380,50){13}
//: {14}(382,48)(428,48){15}
//: {16}(380,46)(380,-26)(344,-26){17}
wire w7;    //: /sn:0 {0}(194,2)(236,2){1}
wire w34;    //: /sn:0 {0}(580,175)(539,175)(539,102)(449,102){1}
wire w25;    //: /sn:0 {0}(428,107)(370,107)(370,109)(311,109){1}
//: {2}(309,107)(309,85)(323,85){3}
//: {4}(307,109)(257,109){5}
wire w4;    //: /sn:0 {0}(257,-152)(306,-152){1}
//: {2}(310,-152)(575,-152)(575,21)(583,21){3}
//: {4}(308,-150)(308,-134)(323,-134){5}
wire w3;    //: /sn:0 {0}(194,-107)(235,-107){1}
wire w22;    //: /sn:0 {0}(428,53)(308,53)(308,58){1}
//: {2}(306,60)(257,60){3}
//: {4}(308,62)(308,80)(323,80){5}
wire w0;    //: /sn:0 {0}(428,261)(387,261)(387,207){1}
//: {2}(389,205)(428,205){3}
//: {4}(387,203)(387,153){5}
//: {6}(389,151)(428,151){7}
//: {8}(387,149)(387,99){9}
//: {10}(389,97)(428,97){11}
//: {12}(387,95)(387,45){13}
//: {14}(389,43)(428,43){15}
//: {16}(387,41)(387,-3){17}
//: {18}(389,-5)(428,-5){19}
//: {20}(387,-7)(387,-91){21}
//: {22}(389,-93)(428,-93){23}
//: {24}(387,-95)(387,-131)(344,-131){25}
wire w30;    //: /sn:0 {0}(194,212)(236,212){1}
wire w37;    //: /sn:0 {0}(449,48)(568,48)(568,31)(583,31){1}
wire w19;    //: /sn:0 {0}(257,0)(306,0){1}
//: {2}(310,0)(428,0){3}
//: {4}(308,-2)(308,-24)(323,-24){5}
wire w23;    //: /sn:0 {0}(449,212)(565,212)(565,180)(580,180){1}
wire w10;    //: /sn:0 {0}(256,-109)(306,-109){1}
//: {2}(310,-109)(555,-109)(555,165)(580,165){3}
//: {4}(308,-111)(308,-129)(323,-129){5}
wire w24;    //: /sn:0 {0}(194,111)(236,111){1}
wire w31;    //: /sn:0 {0}(428,220)(307,220)(307,212){1}
//: {2}(307,208)(307,187)(322,187){3}
//: {4}(305,210)(257,210){5}
wire w1;    //: /sn:0 {0}(194,-155)(236,-155){1}
wire w8;    //: /sn:0 {0}(449,-90)(568,-90)(568,26)(583,26){1}
wire w17;    //: /sn:0 {0}(428,271)(373,271)(373,217){1}
//: {2}(375,215)(428,215){3}
//: {4}(373,213)(373,163){5}
//: {6}(375,161)(428,161){7}
//: {8}(373,159)(373,83)(344,83){9}
wire w28;    //: /sn:0 {0}(428,166)(309,166){1}
//: {2}(307,164)(307,159)(257,159){3}
//: {4}(307,168)(307,182)(322,182){5}
wire w11;    //: /sn:0 {0}(194,156)(236,156){1}
wire w2;    //: /sn:0 {0}(449,158)(573,158)(573,36)(583,36){1}
wire w15;    //: /sn:0 {0}(194,57)(236,57){1}
wire w5;    //: /sn:0 {0}(194,-51)(236,-51){1}
wire w9;    //: /sn:0 {0}(343,185)(367,185)(367,276)(428,276){1}
wire w40;    //: /sn:0 {0}(449,-2)(546,-2)(546,170)(580,170){1}
//: enddecls

  _GGNBUF #(2) g4 (.I(b1), .Z(w24));   //: @(184,111) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g8 (.I0(w1), .I1(b3), .Z(w4));   //: @(247,-152) /sn:0 /w:[ 1 5 0 ]
  _GGAND3 #(8) g44 (.I0(w0), .I1(w6), .I2(w22), .Z(w37));   //: @(439,48) /sn:0 /w:[ 15 15 0 0 ]
  //: IN g16 (b1) @(78,111) /sn:0 /w:[ 0 ]
  _GGNBUF #(2) g3 (.I(b2), .Z(w7));   //: @(184,2) /sn:0 /w:[ 3 0 ]
  //: joint g47 (w0) @(387, 151) /w:[ 6 8 -1 5 ]
  //: IN g17 (b2) @(75,2) /sn:0 /w:[ 0 ]
  //: joint g26 (b2) @(145, 2) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g2 (.I(a2), .Z(w5));   //: @(184,-51) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g23 (.I0(a0), .I1(w30), .Z(w31));   //: @(247,210) /sn:0 /w:[ 0 1 5 ]
  //: joint g30 (a1) @(156, 57) /w:[ 2 -1 1 4 ]
  //: OUT g39 (g) @(663,172) /sn:0 /w:[ 1 ]
  _GGNBUF #(2) g1 (.I(b3), .Z(w3));   //: @(184,-107) /sn:0 /w:[ 3 0 ]
  //: joint g24 (b3) @(143, -107) /w:[ 2 4 1 -1 ]
  //: joint g29 (b1) @(147, 111) /w:[ 2 4 1 -1 ]
  //: joint g60 (w6) @(380, 210) /w:[ 2 4 -1 1 ]
  //: joint g51 (w0) @(387, -93) /w:[ 22 24 -1 21 ]
  //: IN g18 (b3) @(71,-107) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g10 (.I0(w5), .I1(b2), .Z(w16));   //: @(247,-48) /sn:0 /w:[ 1 5 0 ]
  //: joint g25 (a3) @(151, -155) /w:[ 2 -1 1 4 ]
  _GGOR4 #(10) g65 (.I0(w10), .I1(w40), .I2(w34), .I3(w23), .Z(g));   //: @(591,172) /sn:0 /w:[ 3 1 0 1 0 ]
  _GGOR4 #(10) g64 (.I0(w4), .I1(w8), .I2(w37), .I3(w2), .Z(l));   //: @(594,28) /sn:0 /w:[ 3 1 1 1 0 ]
  //: joint g49 (w0) @(387, 43) /w:[ 14 16 -1 13 ]
  _GGNBUF #(2) g6 (.I(b0), .Z(w30));   //: @(184,212) /sn:0 /w:[ 3 0 ]
  //: joint g50 (w0) @(387, 97) /w:[ 10 12 -1 9 ]
  _GGNBUF #(2) g7 (.I(a1), .Z(w15));   //: @(184,57) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g9 (.I0(a3), .I1(w3), .Z(w10));   //: @(246,-109) /sn:0 /w:[ 5 1 0 ]
  _GGNOR2 #(4) g35 (.I0(w28), .I1(w31), .Z(w9));   //: @(333,185) /sn:0 /w:[ 5 3 0 ]
  //: joint g56 (w25) @(309, 109) /w:[ 1 2 4 -1 ]
  //: joint g58 (w28) @(307, 166) /w:[ 1 2 -1 4 ]
  //: IN g22 (a1) @(78,57) /sn:0 /w:[ 0 ]
  //: joint g31 (b0) @(148, 212) /w:[ 2 4 1 -1 ]
  //: joint g59 (w31) @(307, 210) /w:[ -1 2 4 1 ]
  //: joint g67 (w10) @(308, -109) /w:[ 2 4 1 -1 ]
  //: OUT g41 (l) @(661,28) /sn:0 /w:[ 1 ]
  _GGNOR2 #(4) g33 (.I0(w16), .I1(w19), .Z(w6));   //: @(334,-26) /sn:0 /w:[ 5 5 17 ]
  _GGAND2 #(6) g36 (.I0(w0), .I1(w16), .Z(w8));   //: @(439,-90) /sn:0 /w:[ 23 3 0 ]
  _GGAND2 #(6) g45 (.I0(w0), .I1(w19), .Z(w40));   //: @(439,-2) /sn:0 /w:[ 19 3 0 ]
  //: joint g54 (w6) @(380, 48) /w:[ 14 16 -1 13 ]
  //: OUT g40 (e) @(666,268) /sn:0 /w:[ 1 ]
  _GGAND4 #(10) g42 (.I0(w0), .I1(w6), .I2(w17), .I3(w28), .Z(w2));   //: @(439,158) /sn:0 /w:[ 7 7 7 0 0 ]
  //: joint g52 (w16) @(308, -48) /w:[ -1 2 1 4 ]
  //: joint g66 (w4) @(308, -152) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g12 (.I0(w15), .I1(b1), .Z(w22));   //: @(247,60) /sn:0 /w:[ 1 5 3 ]
  //: joint g28 (a0) @(158, 156) /w:[ 2 -1 4 1 ]
  _GGNOR2 #(4) g34 (.I0(w22), .I1(w25), .Z(w17));   //: @(334,83) /sn:0 /w:[ 5 3 9 ]
  //: joint g46 (w0) @(387, 205) /w:[ 2 4 -1 1 ]
  //: joint g57 (w6) @(380, 102) /w:[ 10 12 -1 9 ]
  //: IN g14 (a0) @(79,156) /sn:0 /w:[ 5 ]
  _GGNBUF #(2) g5 (.I(a0), .Z(w11));   //: @(184,156) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g11 (.I0(a2), .I1(w7), .Z(w19));   //: @(247,0) /sn:0 /w:[ 5 1 0 ]
  //: IN g19 (a2) @(73,-51) /sn:0 /w:[ 0 ]
  //: IN g21 (a3) @(72,-155) /sn:0 /w:[ 0 ]
  //: joint g61 (w17) @(373, 215) /w:[ 2 4 -1 1 ]
  //: IN g20 (b0) @(81,212) /sn:0 /w:[ 0 ]
  _GGNOR2 #(4) g32 (.I0(w4), .I1(w10), .Z(w0));   //: @(334,-131) /sn:0 /w:[ 5 5 25 ]
  //: joint g63 (w17) @(373, 161) /w:[ 6 8 -1 5 ]
  _GGNBUF #(2) g0 (.I(a3), .Z(w1));   //: @(184,-155) /sn:0 /w:[ 3 0 ]
  _GGAND2 #(6) g15 (.I0(w11), .I1(b0), .Z(w28));   //: @(247,159) /sn:0 /w:[ 1 5 3 ]
  _GGAND4 #(10) g38 (.I0(w0), .I1(w6), .I2(w17), .I3(w31), .Z(w23));   //: @(439,212) /sn:0 /w:[ 3 3 3 0 0 ]
  _GGAND3 #(8) g43 (.I0(w0), .I1(w6), .I2(w25), .Z(w34));   //: @(439,102) /sn:0 /w:[ 11 11 0 1 ]
  //: joint g27 (a2) @(154, -51) /w:[ 2 -1 1 4 ]
  //: joint g48 (w0) @(387, -5) /w:[ 18 20 -1 17 ]
  _GGAND4 #(10) g37 (.I0(w0), .I1(w6), .I2(w17), .I3(w9), .Z(e));   //: @(439,268) /sn:0 /w:[ 0 0 0 1 0 ]
  //: joint g62 (w6) @(380, 156) /w:[ 6 8 -1 5 ]
  //: joint g55 (w22) @(308, 60) /w:[ -1 1 2 4 ]
  _GGAND2 #(6) g13 (.I0(a1), .I1(w24), .Z(w25));   //: @(247,109) /sn:0 /w:[ 5 1 5 ]
  //: joint g53 (w19) @(308, 0) /w:[ 2 4 1 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin Comp
module Comp(b, a, et, lt, gt);
//: interface  /sz:(63, 64) /bd:[ Li0>b[7:0](32/64) Li1>a[7:0](16/64) Ro0<lt(48/64) Ro1<gt(32/64) Ro2<et(16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output et;    //: /sn:0 {0}(898,-92)(980,-92)(980,-96)(995,-96){1}
input [7:0] b;    //: /sn:0 {0}(#:254,294)(254,276){1}
//: {2}(254,275)(254,230){3}
//: {4}(254,229)(254,189){5}
//: {6}(254,188)(254,145){7}
//: {8}(254,144)(254,-144){9}
//: {10}(254,-145)(254,-190){11}
//: {12}(254,-191)(254,-231){13}
//: {14}(254,-232)(254,-275){15}
//: {16}(254,-276)(254,-496){17}
output lt;    //: /sn:0 {0}(898,194)(995,194){1}
input [7:0] a;    //: /sn:0 {0}(#:192,300)(192,74){1}
//: {2}(192,73)(192,36){3}
//: {4}(192,35)(192,-7){5}
//: {6}(192,-8)(192,-28)(193,-28)(193,-50){7}
//: {8}(193,-51)(193,-198)(192,-198)(192,-346){9}
//: {10}(192,-347)(192,-384){11}
//: {12}(192,-385)(192,-427){13}
//: {14}(192,-428)(192,-471){15}
//: {16}(192,-472)(192,-498){17}
output gt;    //: /sn:0 {0}(898,-380)(980,-380)(980,-382)(995,-382){1}
wire w16;    //: /sn:0 {0}(196,-7)(385,-7)(385,311)(421,311){1}
wire w13;    //: /sn:0 {0}(258,230)(378,230)(378,548)(421,548){1}
wire w6;    //: /sn:0 {0}(196,-384)(422,-384){1}
wire w7;    //: /sn:0 {0}(196,-346)(422,-346){1}
wire w4;    //: /sn:0 {0}(196,-471)(422,-471){1}
wire w25;    //: /sn:0 {0}(802,106)(862,106)(862,191)(877,191){1}
wire w0;    //: /sn:0 {0}(258,-275)(422,-275){1}
wire w3;    //: /sn:0 {0}(258,-144)(422,-144){1}
wire w20;    //: /sn:0 {0}(753,-326)(743,-326)(743,-311)(772,-311)(772,338)(573,338){1}
wire w18;    //: /sn:0 {0}(196,74)(469,74)(469,87){1}
//: {2}(467,89)(461,89){3}
//: {4}(469,91)(469,101)(411,101)(411,392)(421,392){5}
wire w12;    //: /sn:0 {0}(467,204)(472,204){1}
//: {2}(474,202)(474,189)(258,189){3}
//: {4}(474,206)(474,216)(413,216)(413,507)(421,507){5}
wire w19;    //: /sn:0 {0}(781,108)(771,108)(771,123)(790,123)(790,672)(620,672)(620,513)(590,513)(590,501)(573,501){1}
wire w10;    //: /sn:0 {0}(877,-95)(776,-95){1}
//: {2}(772,-95)(661,-95)(661,-328){3}
//: {4}(663,-330)(673,-330)(673,-331)(753,-331){5}
//: {6}(659,-330)(615,-330)(615,-326)(574,-326){7}
//: {8}(774,-93)(774,103)(781,103){9}
wire w23;    //: /sn:0 {0}(774,-328)(862,-328)(862,-378)(877,-378){1}
wire w21;    //: /sn:0 {0}(877,-90)(867,-90)(867,-75)(899,-75)(899,511)(613,511)(613,412)(573,412){1}
wire w1;    //: /sn:0 {0}(258,-231)(422,-231){1}
wire w8;    //: /sn:0 {0}(877,196)(699,196)(699,-237)(574,-237){1}
wire w17;    //: /sn:0 {0}(196,36)(400,36)(400,354)(421,354){1}
wire w14;    //: /sn:0 {0}(258,276)(389,276)(389,594)(421,594){1}
wire w11;    //: /sn:0 {0}(258,145)(474,145)(474,158){1}
//: {2}(472,160)(466,160){3}
//: {4}(474,162)(474,172)(413,172)(413,463)(421,463){5}
wire w2;    //: /sn:0 {0}(258,-190)(422,-190){1}
wire w15;    //: /sn:0 {0}(188,-50)(154,-50)(154,267)(421,267){1}
wire w5;    //: /sn:0 {0}(196,-427)(422,-427){1}
wire w9;    //: /sn:0 {0}(574,-400)(860,-400)(860,-383)(877,-383){1}
//: enddecls

  assign w15 = a[3]; //: TAP g8 @(191,-50) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:0
  assign w14 = b[0]; //: TAP g4 @(252,276) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  assign w4 = a[7]; //: TAP g16 @(190,-471) /sn:0 /R:2 /w:[ 0 15 16 ] /ss:1
  //: IN g3 (b) @(254,296) /sn:0 /R:1 /w:[ 0 ]
  //: joint g26 (w10) @(774, -95) /w:[ 1 -1 2 8 ]
  assign w7 = a[4]; //: TAP g17 @(190,-346) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:1
  //: IN g2 (a) @(192,302) /sn:0 /R:1 /w:[ 0 ]
  comp4 g30 (.a0(w18), .a1(w17), .a2(w16), .a3(w15), .b0(w14), .b1(w13), .b2(w12), .b3(w11), .e(w21), .g(w20), .l(w19));   //: @(422, 213) /sz:(150, 410) /sn:0 /p:[ Li0>5 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Li6>5 Li7>5 Ro0<1 Ro1<1 Ro2<1 ]
  _GGAND2 #(6) g23 (.I0(w10), .I1(w20), .Z(w23));   //: @(764,-328) /sn:0 /w:[ 5 0 0 ]
  //: joint g1 (w18) @(469, 89) /w:[ -1 1 2 4 ]
  _GGAND2 #(6) g24 (.I0(w10), .I1(w19), .Z(w25));   //: @(792,106) /sn:0 /w:[ 9 0 0 ]
  //: OUT g29 (et) @(992,-96) /sn:0 /w:[ 1 ]
  assign w6 = a[5]; //: TAP g18 @(190,-384) /sn:0 /R:2 /w:[ 0 11 12 ] /ss:1
  //: joint g25 (w10) @(661, -330) /w:[ 4 -1 6 3 ]
  assign w17 = a[1]; //: TAP g10 @(190,36) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  assign w12 = b[2]; //: TAP g6 @(252,189) /sn:0 /R:2 /w:[ 3 5 6 ] /ss:1
  assign w16 = a[2]; //: TAP g9 @(190,-7) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:1
  assign w11 = b[3]; //: TAP g7 @(252,145) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  //: joint g31 (w11) @(474, 160) /w:[ -1 1 2 4 ]
  _GGAND2 #(6) g22 (.I0(w10), .I1(w21), .Z(et));   //: @(888,-92) /sn:0 /w:[ 0 0 0 ]
  assign w0 = b[7]; //: TAP g12 @(252,-275) /sn:0 /R:2 /w:[ 0 15 16 ] /ss:1
  //: OUT g28 (lt) @(992,194) /sn:0 /w:[ 1 ]
  assign w2 = b[5]; //: TAP g14 @(252,-190) /sn:0 /R:2 /w:[ 0 11 12 ] /ss:1
  assign w18 = a[0]; //: TAP g11 @(190,74) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  assign w13 = b[1]; //: TAP g5 @(252,230) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  _GGOR2 #(6) g21 (.I0(w25), .I1(w8), .Z(lt));   //: @(888,194) /sn:0 /w:[ 1 0 0 ]
  assign w5 = a[6]; //: TAP g19 @(190,-427) /sn:0 /R:2 /w:[ 0 13 14 ] /ss:1
  //: joint g32 (w12) @(474, 204) /w:[ -1 2 1 4 ]
  _GGOR2 #(6) g20 (.I0(w9), .I1(w23), .Z(gt));   //: @(888,-380) /sn:0 /w:[ 1 1 0 ]
  assign w1 = b[6]; //: TAP g15 @(252,-231) /sn:0 /R:2 /w:[ 0 13 14 ] /ss:1
  comp4 g0 (.a0(w7), .a1(w6), .a2(w5), .a3(w4), .b0(w3), .b1(w2), .b2(w1), .b3(w0), .e(w10), .g(w9), .l(w8));   //: @(423, -525) /sz:(150, 410) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Li6>1 Li7>1 Ro0<7 Ro1<0 Ro2<1 ]
  //: OUT g27 (gt) @(992,-382) /sn:0 /w:[ 1 ]
  assign w3 = b[4]; //: TAP g13 @(252,-144) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin Comparator
module Comparator(B, A, O);
//: interface  /sz:(87, 48) /bd:[ Li0>B[7:0](32/48) Li1>A[7:0](16/48) Ro0<O(16/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:374,49)(453,49){1}
//: {2}(454,49)(472,49){3}
//: {4}(473,49)(493,49){5}
//: {6}(494,49)(514,49){7}
//: {8}(515,49)(533,49){9}
//: {10}(534,49)(553,49){11}
//: {12}(554,49)(569,49){13}
//: {14}(570,49)(588,49){15}
//: {16}(589,49)(609,49){17}
input [7:0] A;    //: /sn:0 {0}(#:83,47)(166,47){1}
//: {2}(167,47)(185,47){3}
//: {4}(186,47)(206,47){5}
//: {6}(207,47)(227,47){7}
//: {8}(228,47)(246,47){9}
//: {10}(247,47)(266,47){11}
//: {12}(267,47)(282,47){13}
//: {14}(283,47)(301,47){15}
//: {16}(302,47)(330,47){17}
output O;    //: /sn:0 {0}(791,313)(812,313)(812,313)(821,313){1}
wire w6;    //: /sn:0 {0}(247,51)(247,338)(648,338){1}
wire w13;    //: /sn:0 {0}(494,53)(494,279)(648,279){1}
wire w16;    //: /sn:0 {0}(473,53)(473,248)(649,248){1}
wire w7;    //: /sn:0 {0}(454,53)(454,217)(644,217){1}
wire w4;    //: /sn:0 {0}(207,51)(207,274)(648,274){1}
wire w39;    //: /sn:0 {0}(770,296)(748,296)(748,215)(665,215){1}
wire w3;    //: /sn:0 {0}(186,51)(186,243)(649,243){1}
wire w36;    //: /sn:0 {0}(770,331)(737,331)(737,409)(669,409){1}
wire w30;    //: /sn:0 {0}(770,321)(726,321)(726,365)(669,365){1}
wire w12;    //: /sn:0 {0}(589,53)(589,411)(648,411){1}
wire w18;    //: /sn:0 {0}(670,246)(741,246)(741,301)(770,301){1}
wire w10;    //: /sn:0 {0}(534,53)(534,343)(648,343){1}
wire w21;    //: /sn:0 {0}(669,277)(735,277)(735,306)(770,306){1}
wire w24;    //: /sn:0 {0}(668,304)(729,304)(729,311)(770,311){1}
wire w1;    //: /sn:0 {0}(267,51)(267,362)(648,362){1}
wire w8;    //: /sn:0 {0}(283,51)(283,384)(648,384){1}
wire w27;    //: /sn:0 {0}(669,341)(722,341)(722,316)(770,316){1}
wire w33;    //: /sn:0 {0}(669,387)(731,387)(731,326)(770,326){1}
wire w14;    //: /sn:0 {0}(515,53)(515,306)(647,306){1}
wire w2;    //: /sn:0 {0}(167,51)(167,212)(644,212){1}
wire w11;    //: /sn:0 {0}(570,53)(570,389)(648,389){1}
wire w15;    //: /sn:0 {0}(554,53)(554,367)(648,367){1}
wire w5;    //: /sn:0 {0}(228,51)(228,301)(647,301){1}
wire w9;    //: /sn:0 {0}(302,51)(302,406)(648,406){1}
//: enddecls

  assign w2 = A[0]; //: TAP g4 @(167,45) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w6 = A[4]; //: TAP g8 @(247,45) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  assign w10 = B[4]; //: TAP g3 @(534,47) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  assign w16 = B[1]; //: TAP g16 @(473,47) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: IN g17 (B) @(372,49) /sn:0 /w:[ 0 ]
  _GGAND8 #(18) g26 (.I0(w39), .I1(w18), .I2(w21), .I3(w24), .I4(w27), .I5(w30), .I6(w33), .I7(w36), .Z(O));   //: @(781,313) /sn:0 /w:[ 0 1 1 1 1 0 1 0 0 ]
  assign w7 = B[0]; //: TAP g2 @(454,47) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  _GGNXOR2 #(6) g23 (.I0(w8), .I1(w11), .Z(w33));   //: @(659,387) /sn:0 /w:[ 1 1 0 ]
  assign w8 = A[6]; //: TAP g1 @(283,45) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  _GGNXOR2 #(6) g24 (.I0(w9), .I1(w12), .Z(w36));   //: @(659,409) /sn:0 /w:[ 1 1 1 ]
  _GGNXOR2 #(6) g18 (.I0(w3), .I1(w16), .Z(w18));   //: @(660,246) /sn:0 /w:[ 1 1 0 ]
  assign w9 = A[7]; //: TAP g10 @(302,45) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  _GGNXOR2 #(6) g25 (.I0(w2), .I1(w7), .Z(w39));   //: @(655,215) /sn:0 /w:[ 1 1 1 ]
  assign w4 = A[2]; //: TAP g6 @(207,45) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w5 = A[3]; //: TAP g7 @(228,45) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w1 = A[5]; //: TAP g9 @(267,45) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  _GGNXOR2 #(6) g22 (.I0(w1), .I1(w15), .Z(w30));   //: @(659,365) /sn:0 /w:[ 1 1 1 ]
  assign w12 = B[7]; //: TAP g12 @(589,47) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  assign w3 = A[1]; //: TAP g5 @(186,45) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign w11 = B[6]; //: TAP g11 @(570,47) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  assign w14 = B[3]; //: TAP g14 @(515,47) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  _GGNXOR2 #(6) g19 (.I0(w4), .I1(w13), .Z(w21));   //: @(659,277) /sn:0 /w:[ 1 1 0 ]
  _GGNXOR2 #(6) g21 (.I0(w6), .I1(w10), .Z(w27));   //: @(659,341) /sn:0 /w:[ 1 1 0 ]
  _GGNXOR2 #(6) g20 (.I0(w5), .I1(w14), .Z(w24));   //: @(658,304) /sn:0 /w:[ 1 1 0 ]
  //: IN g0 (A) @(81,47) /sn:0 /w:[ 0 ]
  assign w15 = B[5]; //: TAP g15 @(554,47) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  //: OUT g27 (O) @(818,313) /sn:0 /w:[ 1 ]
  assign w13 = B[2]; //: TAP g13 @(494,47) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1

endmodule
//: /netlistEnd

